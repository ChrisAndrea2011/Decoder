`ifndef _bp_
`define _bp_
class basepacket;
rand bit enable;
randc bit [3:0] A;
 bit [15:0] Y;
endclass
`endif

